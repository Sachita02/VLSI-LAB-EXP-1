module ha(a,b,sum,carry);
input a,b;
output sum,carry;

module ha (a,b,s,c); 
input a,b; 
output s,c; 
xor g1(s,a,b); 
and g2 (c,a,b); 
endmodule
